// megafunction wizard: %LPM_MUX%VBB%
// GENERATION: STANDARD
// VERSION: WM1.0
// MODULE: lpm_mux 

// ============================================================
// File Name: lpm_mux0.v
// Megafunction Name(s):
// 			lpm_mux
//
// Simulation Library Files(s):
// 			lpm
// ============================================================
// ************************************************************
// THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
//
// 9.1 Build 222 10/21/2009 SJ Web Edition
// ************************************************************

//Copyright (C) 1991-2009 Altera Corporation
//Your use of Altera Corporation's design tools, logic functions 
//and other software and tools, and its AMPP partner logic 
//functions, and any output files from any of the foregoing 
//(including device programming or simulation files), and any 
//associated documentation or information are expressly subject 
//to the terms and conditions of the Altera Program License 
//Subscription Agreement, Altera MegaCore Function License 
//Agreement, or other applicable license agreement, including, 
//without limitation, that your use is for the sole purpose of 
//programming logic devices manufactured by Altera and sold by 
//Altera or its authorized distributors.  Please refer to the 
//applicable agreement for further details.

module lpm_mux0 (
	clken,
	clock,
	data0x,
	data1x,
	data2x,
	data3x,
	data4x,
	data5x,
	data6x,
	data7x,
	sel,
	result);

	input	  clken;
	input	  clock;
	input	[11:0]  data0x;
	input	[11:0]  data1x;
	input	[11:0]  data2x;
	input	[11:0]  data3x;
	input	[11:0]  data4x;
	input	[11:0]  data5x;
	input	[11:0]  data6x;
	input	[11:0]  data7x;
	input	[2:0]  sel;
	output	[11:0]  result;
`ifndef ALTERA_RESERVED_QIS
// synopsys translate_off
`endif
	tri1	  clken;
`ifndef ALTERA_RESERVED_QIS
// synopsys translate_on
`endif

endmodule

// ============================================================
// CNX file retrieval info
// ============================================================
// Retrieval info: PRIVATE: INTENDED_DEVICE_FAMILY STRING "Stratix II"
// Retrieval info: PRIVATE: SYNTH_WRAPPER_GEN_POSTFIX STRING "0"
// Retrieval info: CONSTANT: LPM_PIPELINE NUMERIC "1"
// Retrieval info: CONSTANT: LPM_SIZE NUMERIC "8"
// Retrieval info: CONSTANT: LPM_TYPE STRING "LPM_MUX"
// Retrieval info: CONSTANT: LPM_WIDTH NUMERIC "12"
// Retrieval info: CONSTANT: LPM_WIDTHS NUMERIC "3"
// Retrieval info: USED_PORT: clken 0 0 0 0 INPUT VCC clken
// Retrieval info: USED_PORT: clock 0 0 0 0 INPUT NODEFVAL clock
// Retrieval info: USED_PORT: data0x 0 0 12 0 INPUT NODEFVAL data0x[11..0]
// Retrieval info: USED_PORT: data1x 0 0 12 0 INPUT NODEFVAL data1x[11..0]
// Retrieval info: USED_PORT: data2x 0 0 12 0 INPUT NODEFVAL data2x[11..0]
// Retrieval info: USED_PORT: data3x 0 0 12 0 INPUT NODEFVAL data3x[11..0]
// Retrieval info: USED_PORT: data4x 0 0 12 0 INPUT NODEFVAL data4x[11..0]
// Retrieval info: USED_PORT: data5x 0 0 12 0 INPUT NODEFVAL data5x[11..0]
// Retrieval info: USED_PORT: data6x 0 0 12 0 INPUT NODEFVAL data6x[11..0]
// Retrieval info: USED_PORT: data7x 0 0 12 0 INPUT NODEFVAL data7x[11..0]
// Retrieval info: USED_PORT: result 0 0 12 0 OUTPUT NODEFVAL result[11..0]
// Retrieval info: USED_PORT: sel 0 0 3 0 INPUT NODEFVAL sel[2..0]
// Retrieval info: CONNECT: @clock 0 0 0 0 clock 0 0 0 0
// Retrieval info: CONNECT: @clken 0 0 0 0 clken 0 0 0 0
// Retrieval info: CONNECT: result 0 0 12 0 @result 0 0 12 0
// Retrieval info: CONNECT: @data 0 0 12 84 data7x 0 0 12 0
// Retrieval info: CONNECT: @data 0 0 12 72 data6x 0 0 12 0
// Retrieval info: CONNECT: @data 0 0 12 60 data5x 0 0 12 0
// Retrieval info: CONNECT: @data 0 0 12 48 data4x 0 0 12 0
// Retrieval info: CONNECT: @data 0 0 12 36 data3x 0 0 12 0
// Retrieval info: CONNECT: @data 0 0 12 24 data2x 0 0 12 0
// Retrieval info: CONNECT: @data 0 0 12 12 data1x 0 0 12 0
// Retrieval info: CONNECT: @data 0 0 12 0 data0x 0 0 12 0
// Retrieval info: CONNECT: @sel 0 0 3 0 sel 0 0 3 0
// Retrieval info: LIBRARY: lpm lpm.lpm_components.all
// Retrieval info: GEN_FILE: TYPE_NORMAL lpm_mux0.v TRUE
// Retrieval info: GEN_FILE: TYPE_NORMAL lpm_mux0.inc FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL lpm_mux0.cmp FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL lpm_mux0.bsf TRUE FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL lpm_mux0_inst.v FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL lpm_mux0_bb.v TRUE
// Retrieval info: LIB_FILE: lpm
